`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:05:18 11/09/2010 
// Design Name: 
// Module Name:    indexer32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module indexer32(
	input clk,
	input rst,
	input pse,
	input ld,
	input [31:0] din,
	output dvld,
	output reg [4:0] dout
    );

reg [31:0] match_reg;
wire [31:0] next_match;
reg [31:0] match_mask;

assign next_match = (rst == 1'b1) ? 32'h00000000 : (ld == 1'b1) ? din : (pse == 1'b1) ? match_reg : match_reg & match_mask;

always @(posedge clk) begin
	if (rst)
		match_reg <= 32'h00000000;
	else 
		match_reg <= next_match;
end

assign dvld = (rst == 1'b1) ? 1'b0 : (| match_reg);

always @(match_reg) begin
	casez(match_reg)
	32'b????????_????????_????????_???????1: begin  
		match_mask = 32'b11111111_11111111_11111111_11111110;
		dout = 5'h00;
		end
	32'b????????_????????_????????_??????10: begin  
		match_mask = 32'b11111111_11111111_11111111_11111100;
		dout = 5'h01;
		end
	32'b????????_????????_????????_?????100: begin  
		match_mask = 32'b11111111_11111111_11111111_11111000;
		dout = 5'h02;
		end
	32'b????????_????????_????????_????1000: begin  
		match_mask = 32'b11111111_11111111_11111111_11110000;
		dout = 5'h03;
		end
	32'b????????_????????_????????_???10000: begin  
		match_mask = 32'b11111111_11111111_11111111_11100000;
		dout = 5'h04;
		end
	32'b????????_????????_????????_??100000: begin  
		match_mask = 32'b11111111_11111111_11111111_11000000;
		dout = 5'h05;
		end
	32'b????????_????????_????????_?1000000: begin  
		match_mask = 32'b11111111_11111111_11111111_10000000;
		dout = 5'h06;
		end
	32'b????????_????????_????????_10000000: begin  
		match_mask = 32'b11111111_11111111_11111111_00000000;
		dout = 5'h07;
		end
	
	32'b????????_????????_???????1_00000000: begin  
		match_mask = 32'b11111111_11111111_11111110_00000000;
		dout = 5'h08;
		end
	32'b????????_????????_??????10_00000000: begin  
		match_mask = 32'b11111111_11111111_11111100_00000000;
		dout = 5'h09;
		end
	32'b????????_????????_?????100_00000000: begin  
		match_mask = 32'b11111111_11111111_11111000_00000000;
		dout = 5'h0a;
		end
	32'b????????_????????_????1000_00000000: begin  
		match_mask = 32'b11111111_11111111_11110000_00000000;
		dout = 5'h0b;
		end
	32'b????????_????????_???10000_00000000: begin  
		match_mask = 32'b11111111_11111111_11100000_00000000;
		dout = 5'h0c;
		end
	32'b????????_????????_??100000_00000000: begin  
		match_mask = 32'b11111111_11111111_11000000_00000000;
		dout = 5'h0d;
		end
	32'b????????_????????_?1000000_00000000: begin  
		match_mask = 32'b11111111_11111111_10000000_00000000;
		dout = 5'h0e;
		end
	32'b????????_????????_10000000_00000000: begin  
		match_mask = 32'b11111111_11111111_00000000_00000000;
		dout = 5'h0f;
		end
	
	32'b????????_???????1_00000000_00000000: begin  
		match_mask = 32'b11111111_11111110_00000000_00000000;
		dout = 5'h10;
		end
	32'b????????_??????10_00000000_00000000: begin  
		match_mask = 32'b11111111_11111100_00000000_00000000;
		dout = 5'h11;
		end
	32'b????????_?????100_00000000_00000000: begin  
		match_mask = 32'b11111111_11111000_00000000_00000000;
		dout = 5'h12;
		end
	32'b????????_????1000_00000000_00000000: begin  
		match_mask = 32'b11111111_11110000_00000000_00000000;
		dout = 5'h13;
		end
	32'b????????_???10000_00000000_00000000: begin  
		match_mask = 32'b11111111_11100000_00000000_00000000;
		dout = 5'h14;
		end
	32'b????????_??100000_00000000_00000000: begin  
		match_mask = 32'b11111111_11000000_00000000_00000000;
		dout = 5'h15;
		end
	32'b????????_?1000000_00000000_00000000: begin  
		match_mask = 32'b11111111_10000000_00000000_00000000;
		dout = 5'h16;
		end
	32'b????????_10000000_00000000_00000000: begin  
		match_mask = 32'b11111111_00000000_00000000_00000000;
		dout = 5'h17;
		end
	
	32'b???????1_00000000_00000000_00000000: begin  
		match_mask = 32'b11111110_00000000_00000000_00000000;
		dout = 5'h18;
		end
	32'b??????10_00000000_00000000_00000000: begin  
		match_mask = 32'b11111100_00000000_00000000_00000000;
		dout = 5'h19;
		end
	32'b?????100_00000000_00000000_00000000: begin  
		match_mask = 32'b11111000_00000000_00000000_00000000;
		dout = 5'h1a;
		end
	32'b????1000_00000000_00000000_00000000: begin  
		match_mask = 32'b11110000_00000000_00000000_00000000;
		dout = 5'h1b;
		end
	32'b???10000_00000000_00000000_00000000: begin  
		match_mask = 32'b11100000_00000000_00000000_00000000;
		dout = 5'h1c;
		end
	32'b??100000_00000000_00000000_00000000: begin  
		match_mask = 32'b11000000_00000000_00000000_00000000;
		dout = 5'h1d;
		end
	32'b?1000000_00000000_00000000_00000000: begin  
		match_mask = 32'b10000000_00000000_00000000_00000000;
		dout = 5'h1e;
		end
	32'b10000000_00000000_00000000_00000000: begin  
		match_mask = 32'b00000000_00000000_00000000_00000000;
		dout = 5'h1f;
		end
	default: begin  
		match_mask = 32'b00000000_00000000_00000000_00000000;
		dout = 5'h00;
		end
	endcase
end

endmodule
