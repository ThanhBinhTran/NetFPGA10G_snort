module Protocol_SA_DA #(parameter BVSIZE = 256)(
	input wire [71:0] in,
	output wire [BVSIZE-1:0] outp
	);

	wire [BVSIZE-1:0] w;
	
	assign outp = w;
	
bit_TCAM tcam1 (in, 72'h06_00000000_ac1c0b00, 72'hFF_00000000_ffffff00 , w[0]);
	assign w[1] = w[0];
	assign w[6] = w[0];
	assign w[7] = w[0];
	assign w[14] = w[0];
	assign w[15] = w[0];
	assign w[17] = w[0];
	assign w[19] = w[0];
	assign w[21] = w[0];
	assign w[26] = w[0];
	assign w[27] = w[0];
	assign w[29] = w[0];
	assign w[31] = w[0];
	assign w[34] = w[0];
	assign w[36] = w[0];
	assign w[37] = w[0];
	assign w[40] = w[0];
	assign w[42] = w[0];
	assign w[43] = w[0];
	assign w[44] = w[0];
	assign w[46] = w[0];
	assign w[49] = w[0];
	assign w[50] = w[0];
	assign w[54] = w[0];
	assign w[59] = w[0];
	assign w[61] = w[0];
	assign w[62] = w[0];
	assign w[63] = w[0];
	assign w[68] = w[0];
	assign w[72] = w[0];
	assign w[77] = w[0];
	assign w[83] = w[0];
	assign w[85] = w[0];
	assign w[93] = w[0];
	assign w[94] = w[0];
	assign w[96] = w[0];
	assign w[105] = w[0];
	assign w[119] = w[0];
	assign w[121] = w[0];
	assign w[126] = w[0];
	assign w[133] = w[0];
	assign w[134] = w[0];
	assign w[147] = w[0];
	assign w[158] = w[0];
	assign w[159] = w[0];
	assign w[160] = w[0];
	assign w[162] = w[0];
	assign w[163] = w[0];
	assign w[164] = w[0];
	assign w[165] = w[0];
	assign w[166] = w[0];
	assign w[167] = w[0];
	assign w[170] = w[0];
	assign w[180] = w[0];
	assign w[191] = w[0];
	assign w[193] = w[0];
bit_TCAM tcam2 (in, 72'h06_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[2]);
	assign w[3] = w[2];
	assign w[5] = w[2];
	assign w[8] = w[2];
	assign w[10] = w[2];
	assign w[12] = w[2];
	assign w[20] = w[2];
	assign w[22] = w[2];
	assign w[28] = w[2];
	assign w[30] = w[2];
	assign w[32] = w[2];
	assign w[35] = w[2];
	assign w[39] = w[2];
	assign w[45] = w[2];
	assign w[51] = w[2];
	assign w[52] = w[2];
	assign w[53] = w[2];
	assign w[56] = w[2];
	assign w[57] = w[2];
	assign w[58] = w[2];
	assign w[60] = w[2];
	assign w[65] = w[2];
	assign w[66] = w[2];
	assign w[67] = w[2];
	assign w[69] = w[2];
	assign w[70] = w[2];
	assign w[74] = w[2];
	assign w[75] = w[2];
	assign w[76] = w[2];
	assign w[78] = w[2];
	assign w[79] = w[2];
	assign w[80] = w[2];
	assign w[81] = w[2];
	assign w[82] = w[2];
	assign w[88] = w[2];
	assign w[89] = w[2];
	assign w[90] = w[2];
	assign w[91] = w[2];
	assign w[95] = w[2];
	assign w[98] = w[2];
	assign w[99] = w[2];
	assign w[100] = w[2];
	assign w[101] = w[2];
	assign w[102] = w[2];
	assign w[106] = w[2];
	assign w[107] = w[2];
	assign w[108] = w[2];
	assign w[109] = w[2];
	assign w[110] = w[2];
	assign w[111] = w[2];
	assign w[112] = w[2];
	assign w[113] = w[2];
	assign w[114] = w[2];
	assign w[115] = w[2];
	assign w[116] = w[2];
	assign w[117] = w[2];
	assign w[118] = w[2];
	assign w[120] = w[2];
	assign w[122] = w[2];
	assign w[123] = w[2];
	assign w[124] = w[2];
	assign w[125] = w[2];
	assign w[128] = w[2];
	assign w[129] = w[2];
	assign w[130] = w[2];
	assign w[131] = w[2];
	assign w[135] = w[2];
	assign w[136] = w[2];
	assign w[137] = w[2];
	assign w[138] = w[2];
	assign w[139] = w[2];
	assign w[140] = w[2];
	assign w[141] = w[2];
	assign w[142] = w[2];
	assign w[143] = w[2];
	assign w[144] = w[2];
	assign w[145] = w[2];
	assign w[146] = w[2];
	assign w[150] = w[2];
	assign w[151] = w[2];
	assign w[152] = w[2];
	assign w[153] = w[2];
	assign w[154] = w[2];
	assign w[155] = w[2];
	assign w[156] = w[2];
	assign w[157] = w[2];
	assign w[161] = w[2];
	assign w[168] = w[2];
	assign w[169] = w[2];
	assign w[171] = w[2];
	assign w[172] = w[2];
	assign w[173] = w[2];
	assign w[174] = w[2];
	assign w[175] = w[2];
	assign w[176] = w[2];
	assign w[178] = w[2];
	assign w[179] = w[2];
	assign w[181] = w[2];
	assign w[184] = w[2];
	assign w[185] = w[2];
	assign w[187] = w[2];
	assign w[188] = w[2];
	assign w[189] = w[2];
	assign w[190] = w[2];
	assign w[192] = w[2];
bit_TCAM tcam3 (in, 72'h11_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[4]);
	assign w[23] = w[4];
	assign w[41] = w[4];
	assign w[48] = w[4];
	assign w[55] = w[4];
	assign w[71] = w[4];
	assign w[87] = w[4];
	assign w[182] = w[4];
	assign w[183] = w[4];
	assign w[186] = w[4];
bit_TCAM tcam4 (in, 72'h01_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[9]);
bit_TCAM tcam5 (in, 72'h11_00000000_ac1c0b00, 72'hFF_00000000_ffffff00 , w[11]);
	assign w[25] = w[11];
	assign w[47] = w[11];
	assign w[64] = w[11];
	assign w[73] = w[11];
	assign w[84] = w[11];
	assign w[86] = w[11];
	assign w[92] = w[11];
	assign w[97] = w[11];
	assign w[132] = w[11];
bit_TCAM tcam6 (in, 72'h04_00000000_ac1c0b00, 72'hFF_00000000_ffffff00 , w[13]);
bit_TCAM tcam7 (in, 72'h06_00000000_00000000, 72'hFF_00000000_00000000 , w[16]);
	assign w[18] = w[16];
bit_TCAM tcam8 (in, 72'h11_ac1c0b00_e00000fb, 72'hFF_ffffff00_e00000fb , w[24]);
bit_TCAM tcam9 (in, 72'h01_00000000_ac1c0b00, 72'hFF_00000000_ffffff00 , w[33]);
bit_TCAM tcam10 (in, 72'h06_00000000_00000000, 72'hFF_00000000_00000000 , w[38]);
bit_TCAM tcam11 (in, 72'h06_00000000_00000000, 72'hFF_00000000_00000000 , w[103]);
bit_TCAM tcam12 (in, 72'h11_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[104]);
bit_TCAM tcam13 (in, 72'h06_00000000_00000000, 72'hFF_00000000_00000000 , w[127]);
bit_TCAM tcam14 (in, 72'h06_ac1c0b00_551103fa, 72'hFF_ffffff00_551103fa , w[148]);
bit_TCAM tcam15 (in, 72'h06_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[149]);
bit_TCAM tcam16 (in, 72'h06_ac1c0b00_00000000, 72'hFF_ffffff00_00000000 , w[177]);
bit_TCAM tcam17 (in, 72'h06_00000000_00000000, 72'hFF_00000000_00000000 , w[194]);

endmodule
