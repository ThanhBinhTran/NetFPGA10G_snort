module Group_0(out,clk,sod,eod,en,char,rst);
	input clk, sod, en, eod,rst;
	input [7:0] char;
	output [96:0] out;
	wire [132:0] q_out;

//Centranlized block declare 
	CentralizedCharacter_0 ram (
		.sod(sod),
		.eod(eod),
		.i_char(char),
		.clk(clk),
		.o_match(q_out),
		.en(en));
//Finish centranlized block declare 

//Pcre Engine declare 
	engine_0_0 engine_0_0(
		.out(out[0]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_2(q_out[2]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		.en(en));
	engine_0_1 engine_0_1(
		.out(out[1]), 
		.clk(clk), 
		.sod(sod), 
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_11(q_out[11]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_0(q_out[0]),
		.en(en));
	engine_0_2 engine_0_2(
		.out(out[2]), 
		.clk(clk), 
		.sod(sod), 
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		.en(en));
	engine_0_3 engine_0_3(
		.out(out[3]), 
		.clk(clk), 
		.sod(sod), 
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_23(q_out[23]),
		 .in_1(q_out[1]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_20(q_out[20]),
		.en(en));
	/*
	engine_0_4 engine_0_4(
		.out(out[4]), 
		.clk(clk), 
		.sod(sod), 
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_26(q_out[26]),
		 .in_27(q_out[27]),
		 .in_28(q_out[28]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_31(q_out[31]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		.en(en));
	engine_0_5 engine_0_5(
		.out(out[5]), 
		.clk(clk), 
		.sod(sod), 
		 .in_32(q_out[32]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_27(q_out[27]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_6 engine_0_6(
		.out(out[6]), 
		.clk(clk), 
		.sod(sod), 
		 .in_33(q_out[33]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_26(q_out[26]),
		 .in_27(q_out[27]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_7 engine_0_7(
		.out(out[7]), 
		.clk(clk), 
		.sod(sod), 
		 .in_34(q_out[34]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_8 engine_0_8(
		.out(out[8]), 
		.clk(clk), 
		.sod(sod), 
		 .in_35(q_out[35]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_12(q_out[12]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_9 engine_0_9(
		.out(out[9]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_21(q_out[21]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_27(q_out[27]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_10 engine_0_10(
		.out(out[10]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_12(q_out[12]),
		 .in_21(q_out[21]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_31(q_out[31]),
		.en(en));
	engine_0_11 engine_0_11(
		.out(out[11]), 
		.clk(clk), 
		.sod(sod), 
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_38(q_out[38]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_20(q_out[20]),
		 .in_26(q_out[26]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		.en(en));
	engine_0_12 engine_0_12(
		.out(out[12]), 
		.clk(clk), 
		.sod(sod), 
		 .in_39(q_out[39]),
		 .in_40(q_out[40]),
		 .in_0(q_out[0]),
		 .in_5(q_out[5]),
		 .in_8(q_out[8]),
		 .in_13(q_out[13]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		.en(en));
	engine_0_13 engine_0_13(
		.out(out[13]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_13(q_out[13]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_29(q_out[29]),
		 .in_38(q_out[38]),
		.en(en));
	engine_0_14 engine_0_14(
		.out(out[14]), 
		.clk(clk), 
		.sod(sod), 
		 .in_41(q_out[41]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		.en(en));
	engine_0_15 engine_0_15(
		.out(out[15]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_13(q_out[13]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_16 engine_0_16(
		.out(out[16]), 
		.clk(clk), 
		.sod(sod), 
		 .in_42(q_out[42]),
		 .in_43(q_out[43]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_30(q_out[30]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_17 engine_0_17(
		.out(out[17]), 
		.clk(clk), 
		.sod(sod), 
		 .in_44(q_out[44]),
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		.en(en));
	engine_0_18 engine_0_18(
		.out(out[18]), 
		.clk(clk), 
		.sod(sod), 
		 .in_45(q_out[45]),
		 .in_0(q_out[0]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_14(q_out[14]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_19 engine_0_19(
		.out(out[19]), 
		.clk(clk), 
		.sod(sod), 
		 .in_46(q_out[46]),
		 .in_47(q_out[47]),
		 .in_48(q_out[48]),
		 .in_49(q_out[49]),
		 .in_50(q_out[50]),
		 .in_51(q_out[51]),
		 .in_52(q_out[52]),
		 .in_53(q_out[53]),
		 .in_54(q_out[54]),
		 .in_1(q_out[1]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		.en(en));
	engine_0_20 engine_0_20(
		.out(out[20]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_21 engine_0_21(
		.out(out[21]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_22 engine_0_22(
		.out(out[22]), 
		.clk(clk), 
		.sod(sod), 
		 .in_55(q_out[55]),
		 .in_56(q_out[56]),
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_25(q_out[25]),
		 .in_31(q_out[31]),
		 .in_38(q_out[38]),
		.en(en));
	engine_0_23 engine_0_23(
		.out(out[23]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_38(q_out[38]),
		.en(en));
	engine_0_24 engine_0_24(
		.out(out[24]), 
		.clk(clk), 
		.sod(sod), 
		 .in_57(q_out[57]),
		 .in_3(q_out[3]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_28(q_out[28]),
		.en(en));
	engine_0_25 engine_0_25(
		.out(out[25]), 
		.clk(clk), 
		.sod(sod), 
		 .in_58(q_out[58]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_26 engine_0_26(
		.out(out[26]), 
		.clk(clk), 
		.sod(sod), 
		 .in_59(q_out[59]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_27 engine_0_27(
		.out(out[27]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_26(q_out[26]),
		 .in_37(q_out[37]),
		 .in_45(q_out[45]),
		.en(en));
	engine_0_28 engine_0_28(
		.out(out[28]), 
		.clk(clk), 
		.sod(sod), 
		 .in_60(q_out[60]),
		 .in_61(q_out[61]),
		 .in_62(q_out[62]),
		 .in_63(q_out[63]),
		 .in_64(q_out[64]),
		 .in_65(q_out[65]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_45(q_out[45]),
		 .in_56(q_out[56]),
		.en(en));
	engine_0_29 engine_0_29(
		.out(out[29]), 
		.clk(clk), 
		.sod(sod), 
		 .in_66(q_out[66]),
		 .in_67(q_out[67]),
		 .in_68(q_out[68]),
		 .in_69(q_out[69]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_26(q_out[26]),
		 .in_28(q_out[28]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_58(q_out[58]),
		.en(en));
	engine_0_30 engine_0_30(
		.out(out[30]), 
		.clk(clk), 
		.sod(sod), 
		 .in_70(q_out[70]),
		 .in_71(q_out[71]),
		 .in_72(q_out[72]),
		 .in_73(q_out[73]),
		 .in_74(q_out[74]),
		 .in_75(q_out[75]),
		 .in_76(q_out[76]),
		 .in_77(q_out[77]),
		 .in_78(q_out[78]),
		 .in_79(q_out[79]),
		 .in_80(q_out[80]),
		 .in_81(q_out[81]),
		 .in_13(q_out[13]),
		 .in_20(q_out[20]),
		 .in_33(q_out[33]),
		 .in_49(q_out[49]),
		 .in_51(q_out[51]),
		 .in_57(q_out[57]),
		.en(en));
	engine_0_31 engine_0_31(
		.out(out[31]), 
		.clk(clk), 
		.sod(sod), 
		 .in_82(q_out[82]),
		 .in_83(q_out[83]),
		 .in_84(q_out[84]),
		 .in_85(q_out[85]),
		 .in_86(q_out[86]),
		 .in_87(q_out[87]),
		 .in_88(q_out[88]),
		 .in_89(q_out[89]),
		 .in_90(q_out[90]),
		 .in_91(q_out[91]),
		 .in_1(q_out[1]),
		 .in_25(q_out[25]),
		 .in_46(q_out[46]),
		 .in_51(q_out[51]),
		 .in_57(q_out[57]),
		 .in_75(q_out[75]),
		 .in_79(q_out[79]),
		 .in_81(q_out[81]),
		.en(en));
	engine_0_32 engine_0_32(
		.out(out[32]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_33 engine_0_33(
		.out(out[33]), 
		.clk(clk), 
		.sod(sod), 
		 .in_92(q_out[92]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_22(q_out[22]),
		 .in_30(q_out[30]),
		.en(en));
	engine_0_34 engine_0_34(
		.out(out[34]), 
		.clk(clk), 
		.sod(sod), 
		 .in_93(q_out[93]),
		 .in_94(q_out[94]),
		 .in_95(q_out[95]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_72(q_out[72]),
		 .in_77(q_out[77]),
		.en(en));
	engine_0_35 engine_0_35(
		.out(out[35]), 
		.clk(clk), 
		.sod(sod), 
		 .in_96(q_out[96]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_28(q_out[28]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_57(q_out[57]),
		.en(en));
	engine_0_36 engine_0_36(
		.out(out[36]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_14(q_out[14]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_76(q_out[76]),
		.en(en));
	engine_0_37 engine_0_37(
		.out(out[37]), 
		.clk(clk), 
		.sod(sod), 
		 .in_97(q_out[97]),
		 .in_98(q_out[98]),
		 .in_99(q_out[99]),
		 .in_13(q_out[13]),
		 .in_20(q_out[20]),
		 .in_33(q_out[33]),
		 .in_46(q_out[46]),
		 .in_51(q_out[51]),
		 .in_71(q_out[71]),
		 .in_75(q_out[75]),
		 .in_82(q_out[82]),
		 .in_83(q_out[83]),
		 .in_91(q_out[91]),
		.en(en));
	engine_0_38 engine_0_38(
		.out(out[38]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		.en(en));
	engine_0_39 engine_0_39(
		.out(out[39]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		.en(en));
	engine_0_40 engine_0_40(
		.out(out[40]), 
		.clk(clk), 
		.sod(sod), 
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_19(q_out[19]),
		.en(en));
	engine_0_41 engine_0_41(
		.out(out[41]), 
		.clk(clk), 
		.sod(sod), 
		 .in_102(q_out[102]),
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_56(q_out[56]),
		.en(en));
	engine_0_42 engine_0_42(
		.out(out[42]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_22(q_out[22]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_43 engine_0_43(
		.out(out[43]), 
		.clk(clk), 
		.sod(sod), 
		 .in_2(q_out[2]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_28(q_out[28]),
		 .in_30(q_out[30]),
		 .in_31(q_out[31]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_57(q_out[57]),
		 .in_65(q_out[65]),
		.en(en));
	engine_0_44 engine_0_44(
		.out(out[44]), 
		.clk(clk), 
		.sod(sod), 
		 .in_103(q_out[103]),
		 .in_104(q_out[104]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_20(q_out[20]),
		 .in_28(q_out[28]),
		 .in_57(q_out[57]),
		 .in_74(q_out[74]),
		 .in_78(q_out[78]),
		.en(en));
	engine_0_45 engine_0_45(
		.out(out[45]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_14(q_out[14]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_21(q_out[21]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_44(q_out[44]),
		.en(en));
	engine_0_46 engine_0_46(
		.out(out[46]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_25(q_out[25]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_35(q_out[35]),
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		.en(en));
	engine_0_47 engine_0_47(
		.out(out[47]), 
		.clk(clk), 
		.sod(sod), 
		 .in_105(q_out[105]),
		 .in_0(q_out[0]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_41(q_out[41]),
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		.en(en));
	engine_0_48 engine_0_48(
		.out(out[48]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_2(q_out[2]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_16(q_out[16]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_46(q_out[46]),
		 .in_65(q_out[65]),
		 .in_76(q_out[76]),
		.en(en));
	engine_0_49 engine_0_49(
		.out(out[49]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_37(q_out[37]),
		 .in_56(q_out[56]),
		 .in_63(q_out[63]),
		 .in_65(q_out[65]),
		.en(en));
	engine_0_50 engine_0_50(
		.out(out[50]), 
		.clk(clk), 
		.sod(sod), 
		 .in_106(q_out[106]),
		 .in_107(q_out[107]),
		 .in_108(q_out[108]),
		 .in_1(q_out[1]),
		 .in_31(q_out[31]),
		 .in_33(q_out[33]),
		 .in_46(q_out[46]),
		 .in_50(q_out[50]),
		 .in_70(q_out[70]),
		 .in_72(q_out[72]),
		 .in_74(q_out[74]),
		 .in_77(q_out[77]),
		 .in_79(q_out[79]),
		 .in_83(q_out[83]),
		 .in_87(q_out[87]),
		 .in_90(q_out[90]),
		 .in_97(q_out[97]),
		 .in_99(q_out[99]),
		.en(en));
	engine_0_51 engine_0_51(
		.out(out[51]), 
		.clk(clk), 
		.sod(sod), 
		 .in_109(q_out[109]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		.en(en));
	engine_0_52 engine_0_52(
		.out(out[52]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_43(q_out[43]),
		.en(en));
	engine_0_53 engine_0_53(
		.out(out[53]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_6(q_out[6]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_26(q_out[26]),
		 .in_27(q_out[27]),
		 .in_32(q_out[32]),
		.en(en));
	engine_0_54 engine_0_54(
		.out(out[54]), 
		.clk(clk), 
		.sod(sod), 
		 .in_110(q_out[110]),
		 .in_111(q_out[111]),
		 .in_112(q_out[112]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_20(q_out[20]),
		 .in_22(q_out[22]),
		 .in_26(q_out[26]),
		 .in_30(q_out[30]),
		 .in_39(q_out[39]),
		 .in_41(q_out[41]),
		 .in_42(q_out[42]),
		 .in_44(q_out[44]),
		 .in_55(q_out[55]),
		 .in_57(q_out[57]),
		 .in_98(q_out[98]),
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_55 engine_0_55(
		.out(out[55]), 
		.clk(clk), 
		.sod(sod), 
		 .in_113(q_out[113]),
		 .in_114(q_out[114]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_30(q_out[30]),
		 .in_46(q_out[46]),
		 .in_64(q_out[64]),
		 .in_66(q_out[66]),
		 .in_112(q_out[112]),
		.en(en));
	engine_0_56 engine_0_56(
		.out(out[56]), 
		.clk(clk), 
		.sod(sod), 
		 .in_115(q_out[115]),
		 .in_0(q_out[0]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_25(q_out[25]),
		 .in_30(q_out[30]),
		 .in_31(q_out[31]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_56(q_out[56]),
		 .in_63(q_out[63]),
		 .in_66(q_out[66]),
		.en(en));
	engine_0_57 engine_0_57(
		.out(out[57]), 
		.clk(clk), 
		.sod(sod), 
		 .in_116(q_out[116]),
		 .in_117(q_out[117]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_20(q_out[20]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_101(q_out[101]),
		.en(en));
	engine_0_58 engine_0_58(
		.out(out[58]), 
		.clk(clk), 
		.sod(sod), 
		 .in_118(q_out[118]),
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_69(q_out[69]),
		 .in_105(q_out[105]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_59 engine_0_59(
		.out(out[59]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_110(q_out[110]),
		.en(en));
	engine_0_60 engine_0_60(
		.out(out[60]), 
		.clk(clk), 
		.sod(sod), 
		 .in_119(q_out[119]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_61 engine_0_61(
		.out(out[61]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_119(q_out[119]),
		.en(en));
	engine_0_62 engine_0_62(
		.out(out[62]), 
		.clk(clk), 
		.sod(sod), 
		 .in_120(q_out[120]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_26(q_out[26]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_42(q_out[42]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_63 engine_0_63(
		.out(out[63]), 
		.clk(clk), 
		.sod(sod), 
		 .in_121(q_out[121]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_22(q_out[22]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_42(q_out[42]),
		 .in_43(q_out[43]),
		.en(en));
	engine_0_64 engine_0_64(
		.out(out[64]), 
		.clk(clk), 
		.sod(sod), 
		 .in_122(q_out[122]),
		 .in_123(q_out[123]),
		 .in_124(q_out[124]),
		 .in_125(q_out[125]),
		 .in_4(q_out[4]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_56(q_out[56]),
		 .in_62(q_out[62]),
		 .in_110(q_out[110]),
		.en(en));
	engine_0_65 engine_0_65(
		.out(out[65]), 
		.clk(clk), 
		.sod(sod), 
		 .in_126(q_out[126]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_25(q_out[25]),
		 .in_30(q_out[30]),
		 .in_38(q_out[38]),
		.en(en));
	engine_0_66 engine_0_66(
		.out(out[66]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_22(q_out[22]),
		 .in_25(q_out[25]),
		 .in_26(q_out[26]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_67 engine_0_67(
		.out(out[67]), 
		.clk(clk), 
		.sod(sod), 
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_18(q_out[18]),
		 .in_25(q_out[25]),
		 .in_30(q_out[30]),
		 .in_37(q_out[37]),
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		.en(en));
	engine_0_68 engine_0_68(
		.out(out[68]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_28(q_out[28]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_37(q_out[37]),
		 .in_41(q_out[41]),
		 .in_58(q_out[58]),
		.en(en));
	engine_0_69 engine_0_69(
		.out(out[69]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_26(q_out[26]),
		 .in_28(q_out[28]),
		 .in_29(q_out[29]),
		 .in_32(q_out[32]),
		 .in_35(q_out[35]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_70 engine_0_70(
		.out(out[70]), 
		.clk(clk), 
		.sod(sod), 
		 .in_26(q_out[26]),
		 .in_56(q_out[56]),
		.en(en));
	engine_0_71 engine_0_71(
		.out(out[71]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_20(q_out[20]),
		 .in_21(q_out[21]),
		 .in_24(q_out[24]),
		 .in_25(q_out[25]),
		 .in_28(q_out[28]),
		 .in_56(q_out[56]),
		 .in_57(q_out[57]),
		 .in_65(q_out[65]),
		 .in_66(q_out[66]),
		.en(en));
	engine_0_72 engine_0_72(
		.out(out[72]), 
		.clk(clk), 
		.sod(sod), 
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_20(q_out[20]),
		 .in_25(q_out[25]),
		 .in_28(q_out[28]),
		 .in_35(q_out[35]),
		 .in_60(q_out[60]),
		.en(en));
	engine_0_73 engine_0_73(
		.out(out[73]), 
		.clk(clk), 
		.sod(sod), 
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_12(q_out[12]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_29(q_out[29]),
		 .in_34(q_out[34]),
		 .in_35(q_out[35]),
		.en(en));
	engine_0_74 engine_0_74(
		.out(out[74]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		.en(en));
	engine_0_75 engine_0_75(
		.out(out[75]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_18(q_out[18]),
		 .in_27(q_out[27]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_36(q_out[36]),
		 .in_41(q_out[41]),
		 .in_65(q_out[65]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_76 engine_0_76(
		.out(out[76]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_10(q_out[10]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_35(q_out[35]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		 .in_39(q_out[39]),
		 .in_41(q_out[41]),
		.en(en));
	engine_0_77 engine_0_77(
		.out(out[77]), 
		.clk(clk), 
		.sod(sod), 
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_13(q_out[13]),
		 .in_15(q_out[15]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_29(q_out[29]),
		 .in_35(q_out[35]),
		 .in_46(q_out[46]),
		.en(en));
	engine_0_78 engine_0_78(
		.out(out[78]), 
		.clk(clk), 
		.sod(sod), 
		 .in_127(q_out[127]),
		 .in_12(q_out[12]),
		 .in_28(q_out[28]),
		 .in_78(q_out[78]),
		 .in_81(q_out[81]),
		 .in_90(q_out[90]),
		 .in_94(q_out[94]),
		.en(en));
	engine_0_79 engine_0_79(
		.out(out[79]), 
		.clk(clk), 
		.sod(sod), 
		 .in_2(q_out[2]),
		 .in_5(q_out[5]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_21(q_out[21]),
		 .in_26(q_out[26]),
		 .in_76(q_out[76]),
		.en(en));
	engine_0_80 engine_0_80(
		.out(out[80]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_4(q_out[4]),
		 .in_8(q_out[8]),
		 .in_10(q_out[10]),
		 .in_16(q_out[16]),
		 .in_21(q_out[21]),
		 .in_22(q_out[22]),
		 .in_26(q_out[26]),
		 .in_36(q_out[36]),
		 .in_37(q_out[37]),
		.en(en));
	engine_0_81 engine_0_81(
		.out(out[81]), 
		.clk(clk), 
		.sod(sod), 
		 .in_128(q_out[128]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_41(q_out[41]),
		 .in_76(q_out[76]),
		.en(en));
	engine_0_82 engine_0_82(
		.out(out[82]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_42(q_out[42]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_83 engine_0_83(
		.out(out[83]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_36(q_out[36]),
		 .in_41(q_out[41]),
		 .in_46(q_out[46]),
		.en(en));
	engine_0_84 engine_0_84(
		.out(out[84]), 
		.clk(clk), 
		.sod(sod), 
		 .in_15(q_out[15]),
		 .in_21(q_out[21]),
		 .in_41(q_out[41]),
		 .in_109(q_out[109]),
		.en(en));
	engine_0_85 engine_0_85(
		.out(out[85]), 
		.clk(clk), 
		.sod(sod), 
		 .in_129(q_out[129]),
		 .in_130(q_out[130]),
		 .in_131(q_out[131]),
		 .in_25(q_out[25]),
		 .in_49(q_out[49]),
		 .in_56(q_out[56]),
		 .in_122(q_out[122]),
		.en(en));
	engine_0_86 engine_0_86(
		.out(out[86]), 
		.clk(clk), 
		.sod(sod), 
		 .in_25(q_out[25]),
		 .in_49(q_out[49]),
		 .in_56(q_out[56]),
		 .in_122(q_out[122]),
		 .in_129(q_out[129]),
		 .in_130(q_out[130]),
		 .in_131(q_out[131]),
		.en(en));
	engine_0_87 engine_0_87(
		.out(out[87]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_25(q_out[25]),
		 .in_100(q_out[100]),
		 .in_101(q_out[101]),
		.en(en));
	engine_0_88 engine_0_88(
		.out(out[88]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_29(q_out[29]),
		 .in_30(q_out[30]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_117(q_out[117]),
		.en(en));
	engine_0_89 engine_0_89(
		.out(out[89]), 
		.clk(clk), 
		.sod(sod), 
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_16(q_out[16]),
		 .in_18(q_out[18]),
		 .in_30(q_out[30]),
		 .in_41(q_out[41]),
		 .in_46(q_out[46]),
		.en(en));
	engine_0_90 engine_0_90(
		.out(out[90]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_12(q_out[12]),
		 .in_15(q_out[15]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_20(q_out[20]),
		 .in_32(q_out[32]),
		 .in_42(q_out[42]),
		 .in_65(q_out[65]),
		 .in_110(q_out[110]),
		.en(en));
	engine_0_91 engine_0_91(
		.out(out[91]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_21(q_out[21]),
		 .in_26(q_out[26]),
		.en(en));
	engine_0_92 engine_0_92(
		.out(out[92]), 
		.clk(clk), 
		.sod(sod), 
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_17(q_out[17]),
		 .in_21(q_out[21]),
		 .in_26(q_out[26]),
		 .in_98(q_out[98]),
		 .in_105(q_out[105]),
		.en(en));
	engine_0_93 engine_0_93(
		.out(out[93]), 
		.clk(clk), 
		.sod(sod), 
		 .in_132(q_out[132]),
		 .in_0(q_out[0]),
		 .in_1(q_out[1]),
		 .in_4(q_out[4]),
		 .in_5(q_out[5]),
		 .in_6(q_out[6]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_30(q_out[30]),
		 .in_56(q_out[56]),
		 .in_122(q_out[122]),
		.en(en));
	engine_0_94 engine_0_94(
		.out(out[94]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_6(q_out[6]),
		 .in_7(q_out[7]),
		 .in_8(q_out[8]),
		 .in_9(q_out[9]),
		 .in_12(q_out[12]),
		 .in_14(q_out[14]),
		 .in_15(q_out[15]),
		 .in_16(q_out[16]),
		 .in_17(q_out[17]),
		 .in_18(q_out[18]),
		 .in_19(q_out[19]),
		 .in_26(q_out[26]),
		 .in_27(q_out[27]),
		 .in_30(q_out[30]),
		 .in_32(q_out[32]),
		 .in_35(q_out[35]),
		 .in_38(q_out[38]),
		 .in_41(q_out[41]),
		 .in_42(q_out[42]),
		.en(en));
	engine_0_95 engine_0_95(
		.out(out[95]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_2(q_out[2]),
		 .in_42(q_out[42]),
		 .in_43(q_out[43]),
		.en(en));
	engine_0_96 engine_0_96(
		.out(out[96]), 
		.clk(clk), 
		.sod(sod), 
		 .in_1(q_out[1]),
		 .in_3(q_out[3]),
		 .in_4(q_out[4]),
		 .in_7(q_out[7]),
		 .in_12(q_out[12]),
		 .in_17(q_out[17]),
		 .in_19(q_out[19]),
		 .in_30(q_out[30]),
		 .in_35(q_out[35]),
		 .in_42(q_out[42]),
		.en(en));
*/
//Finish PCRE engine declare 

endmodule
