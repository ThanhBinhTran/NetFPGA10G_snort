module CentralizedCharacter_0(o_match,clk,sod,eod,en,i_char);
	input clk, sod,eod, en;
	input [7:0] i_char;
	output [132:0] o_match;
	wire [132:0] o_ram_0;

	reg [7:0] char_buf;
	//BRAM declare 
	bram_entity_0_0 bram_0 (
		.addr(char_buf),
		.clk(clk),
		.dout(o_ram_0),
		.en(en));
	reg sod_trigger, eod_trigger;
	always@(posedge clk)
	begin
		char_buf <= i_char;
		if(sod)
			sod_trigger <= 1;
		else
			sod_trigger <= 0;
		if(eod)
			eod_trigger <=1;
		else
			eod_trigger <=0;
	end
	assign o_match[0] = sod_trigger | o_ram_0[0];
	assign o_match[1] = o_ram_0[1];
	assign o_match[2] = o_ram_0[2];
	assign o_match[3] = o_ram_0[3];
	assign o_match[4] = o_ram_0[4];
	assign o_match[5] = o_ram_0[5];
	assign o_match[6] = o_ram_0[6];
	assign o_match[7] = o_ram_0[7];
	assign o_match[8] = o_ram_0[8];
	assign o_match[9] = o_ram_0[9];
	assign o_match[10] = o_ram_0[10];
	assign o_match[11] = o_ram_0[11];
	assign o_match[12] = o_ram_0[12];
	assign o_match[13] = o_ram_0[13];
	assign o_match[14] = o_ram_0[14];
	assign o_match[15] = o_ram_0[15];
	assign o_match[16] = o_ram_0[16];
	assign o_match[17] = o_ram_0[17];
	assign o_match[18] = o_ram_0[18];
	assign o_match[19] = o_ram_0[19];
	assign o_match[20] = o_ram_0[20];
	assign o_match[21] = o_ram_0[21];
	assign o_match[22] = o_ram_0[22];
	assign o_match[23] = o_ram_0[23];
	assign o_match[24] = o_ram_0[24];
	assign o_match[25] = o_ram_0[25];
	assign o_match[26] = o_ram_0[26];
	assign o_match[27] = o_ram_0[27];
	assign o_match[28] = o_ram_0[28];
	assign o_match[29] = o_ram_0[29];
	assign o_match[30] = o_ram_0[30];
	assign o_match[31] = o_ram_0[31];
	assign o_match[32] = o_ram_0[32];
	assign o_match[33] = o_ram_0[33];
	assign o_match[34] = o_ram_0[34];
	assign o_match[35] = o_ram_0[35];
	assign o_match[36] = o_ram_0[36];
	assign o_match[37] = o_ram_0[37];
	assign o_match[38] = o_ram_0[38];
	assign o_match[39] = o_ram_0[39];
	assign o_match[40] = o_ram_0[40];
	assign o_match[41] = o_ram_0[41];
	assign o_match[42] = o_ram_0[42];
	assign o_match[43] = o_ram_0[43];
	assign o_match[44] = o_ram_0[44];
	assign o_match[45] = o_ram_0[45];
	assign o_match[46] = sod_trigger | o_ram_0[46];
	assign o_match[47] = o_ram_0[47];
	assign o_match[48] = o_ram_0[48];
	assign o_match[49] = o_ram_0[49];
	assign o_match[50] = o_ram_0[50];
	assign o_match[51] = o_ram_0[51];
	assign o_match[52] = o_ram_0[52];
	assign o_match[53] = o_ram_0[53];
	assign o_match[54] = o_ram_0[54];
	assign o_match[55] = o_ram_0[55];
	assign o_match[56] = o_ram_0[56];
	assign o_match[57] = o_ram_0[57];
	assign o_match[58] = o_ram_0[58];
	assign o_match[59] = o_ram_0[59];
	assign o_match[60] = o_ram_0[60];
	assign o_match[61] = o_ram_0[61];
	assign o_match[62] = o_ram_0[62];
	assign o_match[63] = o_ram_0[63];
	assign o_match[64] = o_ram_0[64];
	assign o_match[65] = o_ram_0[65];
	assign o_match[66] = o_ram_0[66];
	assign o_match[67] = o_ram_0[67];
	assign o_match[68] = o_ram_0[68];
	assign o_match[69] = o_ram_0[69];
	assign o_match[70] = o_ram_0[70];
	assign o_match[71] = o_ram_0[71];
	assign o_match[72] = o_ram_0[72];
	assign o_match[73] = o_ram_0[73];
	assign o_match[74] = o_ram_0[74];
	assign o_match[75] = o_ram_0[75];
	assign o_match[76] = o_ram_0[76];
	assign o_match[77] = o_ram_0[77];
	assign o_match[78] = o_ram_0[78];
	assign o_match[79] = o_ram_0[79];
	assign o_match[80] = o_ram_0[80];
	assign o_match[81] = o_ram_0[81];
	assign o_match[82] = o_ram_0[82];
	assign o_match[83] = o_ram_0[83];
	assign o_match[84] = o_ram_0[84];
	assign o_match[85] = o_ram_0[85];
	assign o_match[86] = o_ram_0[86];
	assign o_match[87] = o_ram_0[87];
	assign o_match[88] = o_ram_0[88];
	assign o_match[89] = o_ram_0[89];
	assign o_match[90] = o_ram_0[90];
	assign o_match[91] = o_ram_0[91];
	assign o_match[92] = o_ram_0[92];
	assign o_match[93] = o_ram_0[93];
	assign o_match[94] = o_ram_0[94];
	assign o_match[95] = o_ram_0[95];
	assign o_match[96] = o_ram_0[96];
	assign o_match[97] = o_ram_0[97];
	assign o_match[98] = o_ram_0[98];
	assign o_match[99] = o_ram_0[99];
	assign o_match[100] = o_ram_0[100];
	assign o_match[101] = o_ram_0[101];
	assign o_match[102] = o_ram_0[102];
	assign o_match[103] = o_ram_0[103];
	assign o_match[104] = o_ram_0[104];
	assign o_match[105] = o_ram_0[105];
	assign o_match[106] = o_ram_0[106];
	assign o_match[107] = o_ram_0[107];
	assign o_match[108] = o_ram_0[108];
	assign o_match[109] = o_ram_0[109];
	assign o_match[110] = o_ram_0[110];
	assign o_match[111] = o_ram_0[111];
	assign o_match[112] = o_ram_0[112];
	assign o_match[113] = o_ram_0[113];
	assign o_match[114] = o_ram_0[114];
	assign o_match[115] = o_ram_0[115];
	assign o_match[116] = o_ram_0[116];
	assign o_match[117] = o_ram_0[117];
	assign o_match[118] = o_ram_0[118];
	assign o_match[119] = o_ram_0[119];
	assign o_match[120] = o_ram_0[120];
	assign o_match[121] = o_ram_0[121];
	assign o_match[122] = o_ram_0[122];
	assign o_match[123] = o_ram_0[123];
	assign o_match[124] = o_ram_0[124];
	assign o_match[125] = o_ram_0[125];
	assign o_match[126] = o_ram_0[126];
	assign o_match[127] = o_ram_0[127];
	assign o_match[128] = o_ram_0[128];
	assign o_match[129] = o_ram_0[129];
	assign o_match[130] = o_ram_0[130];
	assign o_match[131] = o_ram_0[131];
	assign o_match[132] = o_ram_0[132];
endmodule
