module engine_0_38(out,clk,sod,en, in_0, in_1, in_4, in_5, in_8, in_12, in_13, in_15, in_16, in_17, in_18, in_19, in_29, in_30);
//pcre: /^Delta\s+Source\s+\d+\x2E\d+/smi
//block char: ^[9], \x20[8], O[0], L[0], S[0], \x2E[8], \d[5], a[0], r[0], e[0], c[0], d[0], u[0], t[0], 

	input clk,sod,en;

	input in_0, in_1, in_4, in_5, in_8, in_12, in_13, in_15, in_16, in_17, in_18, in_19, in_29, in_30;
	output out;

	assign w0 = 1'b1;
	state_0_38_1 BlockState_0_38_1 (w1,in_0,clk,en,sod,w0);
	state_0_38_2 BlockState_0_38_2 (w2,in_19,clk,en,sod,w1);
	state_0_38_3 BlockState_0_38_3 (w3,in_17,clk,en,sod,w2);
	state_0_38_4 BlockState_0_38_4 (w4,in_5,clk,en,sod,w3);
	state_0_38_5 BlockState_0_38_5 (w5,in_30,clk,en,sod,w4);
	state_0_38_6 BlockState_0_38_6 (w6,in_15,clk,en,sod,w5);
	state_0_38_7 BlockState_0_38_7 (w7,in_1,clk,en,sod,w7,w6);
	state_0_38_8 BlockState_0_38_8 (w8,in_8,clk,en,sod,w7);
	state_0_38_9 BlockState_0_38_9 (w9,in_4,clk,en,sod,w8);
	state_0_38_10 BlockState_0_38_10 (w10,in_29,clk,en,sod,w9);
	state_0_38_11 BlockState_0_38_11 (w11,in_16,clk,en,sod,w10);
	state_0_38_12 BlockState_0_38_12 (w12,in_18,clk,en,sod,w11);
	state_0_38_13 BlockState_0_38_13 (w13,in_17,clk,en,sod,w12);
	state_0_38_14 BlockState_0_38_14 (w14,in_1,clk,en,sod,w14,w13);
	state_0_38_15 BlockState_0_38_15 (w15,in_13,clk,en,sod,w15,w14);
	state_0_38_16 BlockState_0_38_16 (w16,in_12,clk,en,sod,w15);
	state_0_38_17 BlockState_0_38_17 (w17,in_13,clk,en,sod,w17,w16);
	End_state_0_38_18 BlockState_0_38_18 (out,clk,en,sod,w17);
endmodule

module state_0_38_1(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_2(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_3(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_4(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_5(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_6(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_7(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_8(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_9(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_10(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_11(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_12(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_13(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_14(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_15(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_16(out1,in_char,clk,en,rst,in0);
	input in_char,clk,en,rst,in0;
	output out1;
	wire w1,w2;
	assign w1 = in0; 
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module state_0_38_17(out1,in_char,clk,en,rst,in0,in1);
	input in_char,clk,en,rst,in0,in1;
	output out1;
	wire w1,w2;
	or(w1,in0,in1);
	and(w2,in_char,w1);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w2)
);
endmodule

module End_state_0_38_18(out1,clk,en,rst,in0);
	input clk,rst,en,in0;
	output out1;
	wire w1;
	or(w1,out1,in0);
	FDCE #(.INIT(1'b0)) FDCE_inst (
		.Q(out1),
		.C(clk),
		.CE(en),
		.CLR(rst),
		.D(w1)
);
endmodule

